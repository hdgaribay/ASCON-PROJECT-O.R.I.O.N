module constants
	(
	input [3:0] index,
	output reg [63:0] out
	);
	always@(*)begin
		case(index)
			0: out = 64'h00000000000000f0;
			1: out = 64'h00000000000000e1;
			2: out = 64'h00000000000000d2;
			3: out = 64'h00000000000000c3;
			4: out = 64'h00000000000000b4;
			5: out = 64'h00000000000000a5;
			6: out = 64'h0000000000000096;
			7: out = 64'h0000000000000087;
			8: out = 64'h0000000000000078;
			9: out = 64'h0000000000000069;
			10: out = 64'h000000000000005a;
			11: out = 64'h000000000000004b;
			12: out = 64'h000000000000003c;
			13: out = 64'h000000000000002d;
			14: out = 64'h000000000000001e;
			15: out = 64'h000000000000000f;
		endcase
	end
endmodule

